module left_shift_4bit(SllOut, Shift, DataOperand);
    output [31:0] SllOut;
    input Shift;
    input[31:0] DataOperand;
    wire zero;
    assign zero = 0;
    mux2OneBit bit0(SllOut[0], Shift, DataOperand[0], zero);
    mux2OneBit bit1(SllOut[1], Shift, DataOperand[1], zero);
    mux2OneBit bit2(SllOut[2], Shift, DataOperand[2], zero);
    mux2OneBit bit3(SllOut[3], Shift, DataOperand[3], zero);
    mux2OneBit bit4(SllOut[4], Shift, DataOperand[4], zero);
    mux2OneBit bit5(SllOut[5], Shift, DataOperand[5], zero);
    mux2OneBit bit6(SllOut[6], Shift, DataOperand[6], zero);
    mux2OneBit bit7(SllOut[7], Shift, DataOperand[7], zero);
    mux2OneBit bit8(SllOut[8], Shift, DataOperand[8], zero);
    mux2OneBit bit9(SllOut[9], Shift, DataOperand[9], zero);
    mux2OneBit bit10(SllOut[10], Shift, DataOperand[10], zero);
    mux2OneBit bit11(SllOut[11], Shift, DataOperand[11], zero);
    mux2OneBit bit12(SllOut[12], Shift, DataOperand[12], zero);
    mux2OneBit bit13(SllOut[13], Shift, DataOperand[13], zero);
    mux2OneBit bit14(SllOut[14], Shift, DataOperand[14], zero);
    mux2OneBit bit15(SllOut[15], Shift, DataOperand[15], zero);
    mux2OneBit bit16(SllOut[16], Shift, DataOperand[16], DataOperand[0]);
    mux2OneBit bit17(SllOut[17], Shift, DataOperand[17], DataOperand[1]);
    mux2OneBit bit18(SllOut[18], Shift, DataOperand[18], DataOperand[2]);
    mux2OneBit bit19(SllOut[19], Shift, DataOperand[19], DataOperand[3]);
    mux2OneBit bit20(SllOut[20], Shift, DataOperand[20], DataOperand[4]);
    mux2OneBit bit21(SllOut[21], Shift, DataOperand[21], DataOperand[5]);
    mux2OneBit bit22(SllOut[22], Shift, DataOperand[22], DataOperand[6]);
    mux2OneBit bit23(SllOut[23], Shift, DataOperand[23], DataOperand[7]);
    mux2OneBit bit24(SllOut[24], Shift, DataOperand[24], DataOperand[8]);
    mux2OneBit bit25(SllOut[25], Shift, DataOperand[25], DataOperand[9]);
    mux2OneBit bit26(SllOut[26], Shift, DataOperand[26], DataOperand[10]);
    mux2OneBit bit27(SllOut[27], Shift, DataOperand[27], DataOperand[11]);
    mux2OneBit bit28(SllOut[28], Shift, DataOperand[28], DataOperand[12]);
    mux2OneBit bit29(SllOut[29], Shift, DataOperand[29], DataOperand[13]);
    mux2OneBit bit30(SllOut[30], Shift, DataOperand[30], DataOperand[14]);
    mux2OneBit bit31(SllOut[31], Shift, DataOperand[31], DataOperand[15]);
endmodule

module left_shift_3bit(SllOut, Shift, DataOperand);
    output [31:0] SllOut;
    input Shift;
    input[31:0] DataOperand;
    wire zero;
    assign zero = 0;
    mux2OneBit bit0(SllOut[0], Shift, DataOperand[0], zero);
    mux2OneBit bit1(SllOut[1], Shift, DataOperand[1], zero);
    mux2OneBit bit2(SllOut[2], Shift, DataOperand[2], zero);
    mux2OneBit bit3(SllOut[3], Shift, DataOperand[3], zero);
    mux2OneBit bit4(SllOut[4], Shift, DataOperand[4], zero);
    mux2OneBit bit5(SllOut[5], Shift, DataOperand[5], zero);
    mux2OneBit bit6(SllOut[6], Shift, DataOperand[6], zero);
    mux2OneBit bit7(SllOut[7], Shift, DataOperand[7], zero);
    mux2OneBit bit8(SllOut[8], Shift, DataOperand[8], DataOperand[0]);
    mux2OneBit bit9(SllOut[9], Shift, DataOperand[9], DataOperand[1]);
    mux2OneBit bit10(SllOut[10], Shift, DataOperand[10], DataOperand[2]);
    mux2OneBit bit11(SllOut[11], Shift, DataOperand[11], DataOperand[3]);
    mux2OneBit bit12(SllOut[12], Shift, DataOperand[12], DataOperand[4]);
    mux2OneBit bit13(SllOut[13], Shift, DataOperand[13], DataOperand[5]);
    mux2OneBit bit14(SllOut[14], Shift, DataOperand[14], DataOperand[6]);
    mux2OneBit bit15(SllOut[15], Shift, DataOperand[15], DataOperand[7]);
    mux2OneBit bit16(SllOut[16], Shift, DataOperand[16], DataOperand[8]);
    mux2OneBit bit17(SllOut[17], Shift, DataOperand[17], DataOperand[9]);
    mux2OneBit bit18(SllOut[18], Shift, DataOperand[18], DataOperand[10]);
    mux2OneBit bit19(SllOut[19], Shift, DataOperand[19], DataOperand[11]);
    mux2OneBit bit20(SllOut[20], Shift, DataOperand[20], DataOperand[12]);
    mux2OneBit bit21(SllOut[21], Shift, DataOperand[21], DataOperand[13]);
    mux2OneBit bit22(SllOut[22], Shift, DataOperand[22], DataOperand[14]);
    mux2OneBit bit23(SllOut[23], Shift, DataOperand[23], DataOperand[15]);
    mux2OneBit bit24(SllOut[24], Shift, DataOperand[24], DataOperand[16]);
    mux2OneBit bit25(SllOut[25], Shift, DataOperand[25], DataOperand[17]);
    mux2OneBit bit26(SllOut[26], Shift, DataOperand[26], DataOperand[18]);
    mux2OneBit bit27(SllOut[27], Shift, DataOperand[27], DataOperand[19]);
    mux2OneBit bit28(SllOut[28], Shift, DataOperand[28], DataOperand[20]);
    mux2OneBit bit29(SllOut[29], Shift, DataOperand[29], DataOperand[21]);
    mux2OneBit bit30(SllOut[30], Shift, DataOperand[30], DataOperand[22]);
    mux2OneBit bit31(SllOut[31], Shift, DataOperand[31], DataOperand[23]);
endmodule

module left_shift_2bit(SllOut, Shift, DataOperand);
    output [31:0] SllOut;
    input Shift;
    input[31:0] DataOperand;
    wire zero;
    assign zero = 0;
    mux2OneBit bit0(SllOut[0], Shift, DataOperand[0], zero);
    mux2OneBit bit1(SllOut[1], Shift, DataOperand[1], zero);
    mux2OneBit bit2(SllOut[2], Shift, DataOperand[2], zero);
    mux2OneBit bit3(SllOut[3], Shift, DataOperand[3], zero);
    mux2OneBit bit4(SllOut[4], Shift, DataOperand[4], DataOperand[0]);
    mux2OneBit bit5(SllOut[5], Shift, DataOperand[5], DataOperand[1]);
    mux2OneBit bit6(SllOut[6], Shift, DataOperand[6], DataOperand[2]);
    mux2OneBit bit7(SllOut[7], Shift, DataOperand[7], DataOperand[3]);
    mux2OneBit bit8(SllOut[8], Shift, DataOperand[8], DataOperand[4]);
    mux2OneBit bit9(SllOut[9], Shift, DataOperand[9], DataOperand[5]);
    mux2OneBit bit10(SllOut[10], Shift, DataOperand[10], DataOperand[6]);
    mux2OneBit bit11(SllOut[11], Shift, DataOperand[11], DataOperand[7]);
    mux2OneBit bit12(SllOut[12], Shift, DataOperand[12], DataOperand[8]);
    mux2OneBit bit13(SllOut[13], Shift, DataOperand[13], DataOperand[9]);
    mux2OneBit bit14(SllOut[14], Shift, DataOperand[14], DataOperand[10]);
    mux2OneBit bit15(SllOut[15], Shift, DataOperand[15], DataOperand[11]);
    mux2OneBit bit16(SllOut[16], Shift, DataOperand[16], DataOperand[12]);
    mux2OneBit bit17(SllOut[17], Shift, DataOperand[17], DataOperand[13]);
    mux2OneBit bit18(SllOut[18], Shift, DataOperand[18], DataOperand[14]);
    mux2OneBit bit19(SllOut[19], Shift, DataOperand[19], DataOperand[15]);
    mux2OneBit bit20(SllOut[20], Shift, DataOperand[20], DataOperand[16]);
    mux2OneBit bit21(SllOut[21], Shift, DataOperand[21], DataOperand[17]);
    mux2OneBit bit22(SllOut[22], Shift, DataOperand[22], DataOperand[18]);
    mux2OneBit bit23(SllOut[23], Shift, DataOperand[23], DataOperand[19]);
    mux2OneBit bit24(SllOut[24], Shift, DataOperand[24], DataOperand[20]);
    mux2OneBit bit25(SllOut[25], Shift, DataOperand[25], DataOperand[21]);
    mux2OneBit bit26(SllOut[26], Shift, DataOperand[26], DataOperand[22]);
    mux2OneBit bit27(SllOut[27], Shift, DataOperand[27], DataOperand[23]);
    mux2OneBit bit28(SllOut[28], Shift, DataOperand[28], DataOperand[24]);
    mux2OneBit bit29(SllOut[29], Shift, DataOperand[29], DataOperand[25]);
    mux2OneBit bit30(SllOut[30], Shift, DataOperand[30], DataOperand[26]);
    mux2OneBit bit31(SllOut[31], Shift, DataOperand[31], DataOperand[27]);
endmodule

module left_shift_1bit(SllOut, Shift, DataOperand);
    output [31:0] SllOut;
    input Shift;
    input[31:0] DataOperand;
    wire zero;
    assign zero = 0;
    mux2OneBit bit0(SllOut[0], Shift, DataOperand[0], zero);
    mux2OneBit bit1(SllOut[1], Shift, DataOperand[1], zero);
    mux2OneBit bit2(SllOut[2], Shift, DataOperand[2], DataOperand[0]);
    mux2OneBit bit3(SllOut[3], Shift, DataOperand[3], DataOperand[1]);
    mux2OneBit bit4(SllOut[4], Shift, DataOperand[4], DataOperand[2]);
    mux2OneBit bit5(SllOut[5], Shift, DataOperand[5], DataOperand[3]);
    mux2OneBit bit6(SllOut[6], Shift, DataOperand[6], DataOperand[4]);
    mux2OneBit bit7(SllOut[7], Shift, DataOperand[7], DataOperand[5]);
    mux2OneBit bit8(SllOut[8], Shift, DataOperand[8], DataOperand[6]);
    mux2OneBit bit9(SllOut[9], Shift, DataOperand[9], DataOperand[7]);
    mux2OneBit bit10(SllOut[10], Shift, DataOperand[10], DataOperand[8]);
    mux2OneBit bit11(SllOut[11], Shift, DataOperand[11], DataOperand[9]);
    mux2OneBit bit12(SllOut[12], Shift, DataOperand[12], DataOperand[10]);
    mux2OneBit bit13(SllOut[13], Shift, DataOperand[13], DataOperand[11]);
    mux2OneBit bit14(SllOut[14], Shift, DataOperand[14], DataOperand[12]);
    mux2OneBit bit15(SllOut[15], Shift, DataOperand[15], DataOperand[13]);
    mux2OneBit bit16(SllOut[16], Shift, DataOperand[16], DataOperand[14]);
    mux2OneBit bit17(SllOut[17], Shift, DataOperand[17], DataOperand[15]);
    mux2OneBit bit18(SllOut[18], Shift, DataOperand[18], DataOperand[16]);
    mux2OneBit bit19(SllOut[19], Shift, DataOperand[19], DataOperand[17]);
    mux2OneBit bit20(SllOut[20], Shift, DataOperand[20], DataOperand[18]);
    mux2OneBit bit21(SllOut[21], Shift, DataOperand[21], DataOperand[19]);
    mux2OneBit bit22(SllOut[22], Shift, DataOperand[22], DataOperand[20]);
    mux2OneBit bit23(SllOut[23], Shift, DataOperand[23], DataOperand[21]);
    mux2OneBit bit24(SllOut[24], Shift, DataOperand[24], DataOperand[22]);
    mux2OneBit bit25(SllOut[25], Shift, DataOperand[25], DataOperand[23]);
    mux2OneBit bit26(SllOut[26], Shift, DataOperand[26], DataOperand[24]);
    mux2OneBit bit27(SllOut[27], Shift, DataOperand[27], DataOperand[25]);
    mux2OneBit bit28(SllOut[28], Shift, DataOperand[28], DataOperand[26]);
    mux2OneBit bit29(SllOut[29], Shift, DataOperand[29], DataOperand[27]);
    mux2OneBit bit30(SllOut[30], Shift, DataOperand[30], DataOperand[28]);
    mux2OneBit bit31(SllOut[31], Shift, DataOperand[31], DataOperand[29]);
endmodule

module left_shift_0bit(SllOut, Shift, DataOperand);
    output [31:0] SllOut;
    input Shift;
    input[31:0] DataOperand;
    wire zero;
    assign zero = 0;
    mux2OneBit bit0(SllOut[0], Shift, DataOperand[0], zero);
    mux2OneBit bit1(SllOut[1], Shift, DataOperand[1], DataOperand[0]);
    mux2OneBit bit2(SllOut[2], Shift, DataOperand[2], DataOperand[1]);
    mux2OneBit bit3(SllOut[3], Shift, DataOperand[3], DataOperand[2]);
    mux2OneBit bit4(SllOut[4], Shift, DataOperand[4], DataOperand[3]);
    mux2OneBit bit5(SllOut[5], Shift, DataOperand[5], DataOperand[4]);
    mux2OneBit bit6(SllOut[6], Shift, DataOperand[6], DataOperand[5]);
    mux2OneBit bit7(SllOut[7], Shift, DataOperand[7], DataOperand[6]);
    mux2OneBit bit8(SllOut[8], Shift, DataOperand[8], DataOperand[7]);
    mux2OneBit bit9(SllOut[9], Shift, DataOperand[9], DataOperand[8]);
    mux2OneBit bit10(SllOut[10], Shift, DataOperand[10], DataOperand[9]);
    mux2OneBit bit11(SllOut[11], Shift, DataOperand[11], DataOperand[10]);
    mux2OneBit bit12(SllOut[12], Shift, DataOperand[12], DataOperand[11]);
    mux2OneBit bit13(SllOut[13], Shift, DataOperand[13], DataOperand[12]);
    mux2OneBit bit14(SllOut[14], Shift, DataOperand[14], DataOperand[13]);
    mux2OneBit bit15(SllOut[15], Shift, DataOperand[15], DataOperand[14]);
    mux2OneBit bit16(SllOut[16], Shift, DataOperand[16], DataOperand[15]);
    mux2OneBit bit17(SllOut[17], Shift, DataOperand[17], DataOperand[16]);
    mux2OneBit bit18(SllOut[18], Shift, DataOperand[18], DataOperand[17]);
    mux2OneBit bit19(SllOut[19], Shift, DataOperand[19], DataOperand[18]);
    mux2OneBit bit20(SllOut[20], Shift, DataOperand[20], DataOperand[19]);
    mux2OneBit bit21(SllOut[21], Shift, DataOperand[21], DataOperand[20]);
    mux2OneBit bit22(SllOut[22], Shift, DataOperand[22], DataOperand[21]);
    mux2OneBit bit23(SllOut[23], Shift, DataOperand[23], DataOperand[22]);
    mux2OneBit bit24(SllOut[24], Shift, DataOperand[24], DataOperand[23]);
    mux2OneBit bit25(SllOut[25], Shift, DataOperand[25], DataOperand[24]);
    mux2OneBit bit26(SllOut[26], Shift, DataOperand[26], DataOperand[25]);
    mux2OneBit bit27(SllOut[27], Shift, DataOperand[27], DataOperand[26]);
    mux2OneBit bit28(SllOut[28], Shift, DataOperand[28], DataOperand[27]);
    mux2OneBit bit29(SllOut[29], Shift, DataOperand[29], DataOperand[28]);
    mux2OneBit bit30(SllOut[30], Shift, DataOperand[30], DataOperand[29]);
    mux2OneBit bit31(SllOut[31], Shift, DataOperand[31], DataOperand[30]);
endmodule


module left_shifter(SllOut, ShiftAmt, DataOperand);
    input [31:0] DataOperand;
    input[4:0] ShiftAmt;
    output[31:0] SllOut;
    wire [31:0] Bit0Res, Bit1Res, Bit2Res, Bit3Res, Bit4Res;
    left_shift_0bit leftShift0(Bit0Res, ShiftAmt[0], DataOperand);
    left_shift_1bit leftShift1(Bit1Res, ShiftAmt[1], Bit0Res);
    left_shift_2bit leftShift2(Bit2Res, ShiftAmt[2], Bit1Res);
    left_shift_3bit leftShift3(Bit3Res, ShiftAmt[3], Bit2Res);
    left_shift_4bit leftShift4(SllOut, ShiftAmt[4], Bit3Res);
endmodule

module right_shift_4bit(SraOut, Shift, DataOperand);
    output [31:0] SraOut;
    input Shift;
    input[31:0] DataOperand;
    wire ones;
    assign ones = DataOperand[31];
    mux2OneBit bit0(SraOut[0], Shift, DataOperand[0], DataOperand[16]);
    mux2OneBit bit1(SraOut[1], Shift, DataOperand[1], DataOperand[17]);
    mux2OneBit bit2(SraOut[2], Shift, DataOperand[2], DataOperand[18]);
    mux2OneBit bit3(SraOut[3], Shift, DataOperand[3], DataOperand[19]);
    mux2OneBit bit4(SraOut[4], Shift, DataOperand[4], DataOperand[20]);
    mux2OneBit bit5(SraOut[5], Shift, DataOperand[5], DataOperand[21]);
    mux2OneBit bit6(SraOut[6], Shift, DataOperand[6], DataOperand[22]);
    mux2OneBit bit7(SraOut[7], Shift, DataOperand[7], DataOperand[23]);
    mux2OneBit bit8(SraOut[8], Shift, DataOperand[8], DataOperand[24]);
    mux2OneBit bit9(SraOut[9], Shift, DataOperand[9], DataOperand[25]);
    mux2OneBit bit10(SraOut[10], Shift, DataOperand[10], DataOperand[26]);
    mux2OneBit bit11(SraOut[11], Shift, DataOperand[11], DataOperand[27]);
    mux2OneBit bit12(SraOut[12], Shift, DataOperand[12], DataOperand[28]);
    mux2OneBit bit13(SraOut[13], Shift, DataOperand[13], DataOperand[29]);
    mux2OneBit bit14(SraOut[14], Shift, DataOperand[14], DataOperand[30]);
    mux2OneBit bit15(SraOut[15], Shift, DataOperand[15], DataOperand[31]);
    mux2OneBit bit16(SraOut[16], Shift, DataOperand[16], ones);
    mux2OneBit bit17(SraOut[17], Shift, DataOperand[17], ones);
    mux2OneBit bit18(SraOut[18], Shift, DataOperand[18], ones);
    mux2OneBit bit19(SraOut[19], Shift, DataOperand[19], ones);
    mux2OneBit bit20(SraOut[20], Shift, DataOperand[20], ones);
    mux2OneBit bit21(SraOut[21], Shift, DataOperand[21], ones);
    mux2OneBit bit22(SraOut[22], Shift, DataOperand[22], ones);
    mux2OneBit bit23(SraOut[23], Shift, DataOperand[23], ones);
    mux2OneBit bit24(SraOut[24], Shift, DataOperand[24], ones);
    mux2OneBit bit25(SraOut[25], Shift, DataOperand[25], ones);
    mux2OneBit bit26(SraOut[26], Shift, DataOperand[26], ones);
    mux2OneBit bit27(SraOut[27], Shift, DataOperand[27], ones);
    mux2OneBit bit28(SraOut[28], Shift, DataOperand[28], ones);
    mux2OneBit bit29(SraOut[29], Shift, DataOperand[29], ones);
    mux2OneBit bit30(SraOut[30], Shift, DataOperand[30], ones);
    mux2OneBit bit31(SraOut[31], Shift, DataOperand[31], ones);
endmodule

module right_shift_3bit(SraOut, Shift, DataOperand);
    output [31:0] SraOut;
    input Shift;
    input[31:0] DataOperand;
    wire ones;
    assign ones = DataOperand[31];
    mux2OneBit bit0(SraOut[0], Shift, DataOperand[0], DataOperand[8]);
    mux2OneBit bit1(SraOut[1], Shift, DataOperand[1], DataOperand[9]);
    mux2OneBit bit2(SraOut[2], Shift, DataOperand[2], DataOperand[10]);
    mux2OneBit bit3(SraOut[3], Shift, DataOperand[3], DataOperand[11]);
    mux2OneBit bit4(SraOut[4], Shift, DataOperand[4], DataOperand[12]);
    mux2OneBit bit5(SraOut[5], Shift, DataOperand[5], DataOperand[13]);
    mux2OneBit bit6(SraOut[6], Shift, DataOperand[6], DataOperand[14]);
    mux2OneBit bit7(SraOut[7], Shift, DataOperand[7], DataOperand[15]);
    mux2OneBit bit8(SraOut[8], Shift, DataOperand[8], DataOperand[16]);
    mux2OneBit bit9(SraOut[9], Shift, DataOperand[9], DataOperand[17]);
    mux2OneBit bit10(SraOut[10], Shift, DataOperand[10], DataOperand[18]);
    mux2OneBit bit11(SraOut[11], Shift, DataOperand[11], DataOperand[19]);
    mux2OneBit bit12(SraOut[12], Shift, DataOperand[12], DataOperand[20]);
    mux2OneBit bit13(SraOut[13], Shift, DataOperand[13], DataOperand[21]);
    mux2OneBit bit14(SraOut[14], Shift, DataOperand[14], DataOperand[22]);
    mux2OneBit bit15(SraOut[15], Shift, DataOperand[15], DataOperand[23]);
    mux2OneBit bit16(SraOut[16], Shift, DataOperand[16], DataOperand[24]);
    mux2OneBit bit17(SraOut[17], Shift, DataOperand[17], DataOperand[25]);
    mux2OneBit bit18(SraOut[18], Shift, DataOperand[18], DataOperand[26]);
    mux2OneBit bit19(SraOut[19], Shift, DataOperand[19], DataOperand[27]);
    mux2OneBit bit20(SraOut[20], Shift, DataOperand[20], DataOperand[28]);
    mux2OneBit bit21(SraOut[21], Shift, DataOperand[21], DataOperand[29]);
    mux2OneBit bit22(SraOut[22], Shift, DataOperand[22], DataOperand[30]);
    mux2OneBit bit23(SraOut[23], Shift, DataOperand[23], DataOperand[31]);
    mux2OneBit bit24(SraOut[24], Shift, DataOperand[24], ones);
    mux2OneBit bit25(SraOut[25], Shift, DataOperand[25], ones);
    mux2OneBit bit26(SraOut[26], Shift, DataOperand[26], ones);
    mux2OneBit bit27(SraOut[27], Shift, DataOperand[27], ones);
    mux2OneBit bit28(SraOut[28], Shift, DataOperand[28], ones);
    mux2OneBit bit29(SraOut[29], Shift, DataOperand[29], ones);
    mux2OneBit bit30(SraOut[30], Shift, DataOperand[30], ones);
    mux2OneBit bit31(SraOut[31], Shift, DataOperand[31], ones);
endmodule

module right_shift_2bit(SraOut, Shift, DataOperand);
    output [31:0] SraOut;
    input Shift;
    input[31:0] DataOperand;
    wire ones;
    assign ones = DataOperand[31];
    mux2OneBit bit0(SraOut[0], Shift, DataOperand[0], DataOperand[4]);
    mux2OneBit bit1(SraOut[1], Shift, DataOperand[1], DataOperand[5]);
    mux2OneBit bit2(SraOut[2], Shift, DataOperand[2], DataOperand[6]);
    mux2OneBit bit3(SraOut[3], Shift, DataOperand[3], DataOperand[7]);
    mux2OneBit bit4(SraOut[4], Shift, DataOperand[4], DataOperand[8]);
    mux2OneBit bit5(SraOut[5], Shift, DataOperand[5], DataOperand[9]);
    mux2OneBit bit6(SraOut[6], Shift, DataOperand[6], DataOperand[10]);
    mux2OneBit bit7(SraOut[7], Shift, DataOperand[7], DataOperand[11]);
    mux2OneBit bit8(SraOut[8], Shift, DataOperand[8], DataOperand[12]);
    mux2OneBit bit9(SraOut[9], Shift, DataOperand[9], DataOperand[13]);
    mux2OneBit bit10(SraOut[10], Shift, DataOperand[10], DataOperand[14]);
    mux2OneBit bit11(SraOut[11], Shift, DataOperand[11], DataOperand[15]);
    mux2OneBit bit12(SraOut[12], Shift, DataOperand[12], DataOperand[16]);
    mux2OneBit bit13(SraOut[13], Shift, DataOperand[13], DataOperand[17]);
    mux2OneBit bit14(SraOut[14], Shift, DataOperand[14], DataOperand[18]);
    mux2OneBit bit15(SraOut[15], Shift, DataOperand[15], DataOperand[19]);
    mux2OneBit bit16(SraOut[16], Shift, DataOperand[16], DataOperand[20]);
    mux2OneBit bit17(SraOut[17], Shift, DataOperand[17], DataOperand[21]);
    mux2OneBit bit18(SraOut[18], Shift, DataOperand[18], DataOperand[22]);
    mux2OneBit bit19(SraOut[19], Shift, DataOperand[19], DataOperand[23]);
    mux2OneBit bit20(SraOut[20], Shift, DataOperand[20], DataOperand[24]);
    mux2OneBit bit21(SraOut[21], Shift, DataOperand[21], DataOperand[25]);
    mux2OneBit bit22(SraOut[22], Shift, DataOperand[22], DataOperand[26]);
    mux2OneBit bit23(SraOut[23], Shift, DataOperand[23], DataOperand[27]);
    mux2OneBit bit24(SraOut[24], Shift, DataOperand[24], DataOperand[28]);
    mux2OneBit bit25(SraOut[25], Shift, DataOperand[25], DataOperand[29]);
    mux2OneBit bit26(SraOut[26], Shift, DataOperand[26], DataOperand[30]);
    mux2OneBit bit27(SraOut[27], Shift, DataOperand[27], DataOperand[31]);
    mux2OneBit bit28(SraOut[28], Shift, DataOperand[28], ones);
    mux2OneBit bit29(SraOut[29], Shift, DataOperand[29], ones);
    mux2OneBit bit30(SraOut[30], Shift, DataOperand[30], ones);
    mux2OneBit bit31(SraOut[31], Shift, DataOperand[31], ones);
endmodule

module right_shift_1bit(SraOut, Shift, DataOperand);
    output [31:0] SraOut;
    input Shift;
    input[31:0] DataOperand;
    wire ones;
    assign ones = DataOperand[31];
    mux2OneBit bit0(SraOut[0], Shift, DataOperand[0], DataOperand[2]);
    mux2OneBit bit1(SraOut[1], Shift, DataOperand[1], DataOperand[3]);
    mux2OneBit bit2(SraOut[2], Shift, DataOperand[2], DataOperand[4]);
    mux2OneBit bit3(SraOut[3], Shift, DataOperand[3], DataOperand[5]);
    mux2OneBit bit4(SraOut[4], Shift, DataOperand[4], DataOperand[6]);
    mux2OneBit bit5(SraOut[5], Shift, DataOperand[5], DataOperand[7]);
    mux2OneBit bit6(SraOut[6], Shift, DataOperand[6], DataOperand[8]);
    mux2OneBit bit7(SraOut[7], Shift, DataOperand[7], DataOperand[9]);
    mux2OneBit bit8(SraOut[8], Shift, DataOperand[8], DataOperand[10]);
    mux2OneBit bit9(SraOut[9], Shift, DataOperand[9], DataOperand[11]);
    mux2OneBit bit10(SraOut[10], Shift, DataOperand[10], DataOperand[12]);
    mux2OneBit bit11(SraOut[11], Shift, DataOperand[11], DataOperand[13]);
    mux2OneBit bit12(SraOut[12], Shift, DataOperand[12], DataOperand[14]);
    mux2OneBit bit13(SraOut[13], Shift, DataOperand[13], DataOperand[15]);
    mux2OneBit bit14(SraOut[14], Shift, DataOperand[14], DataOperand[16]);
    mux2OneBit bit15(SraOut[15], Shift, DataOperand[15], DataOperand[17]);
    mux2OneBit bit16(SraOut[16], Shift, DataOperand[16], DataOperand[18]);
    mux2OneBit bit17(SraOut[17], Shift, DataOperand[17], DataOperand[19]);
    mux2OneBit bit18(SraOut[18], Shift, DataOperand[18], DataOperand[20]);
    mux2OneBit bit19(SraOut[19], Shift, DataOperand[19], DataOperand[21]);
    mux2OneBit bit20(SraOut[20], Shift, DataOperand[20], DataOperand[22]);
    mux2OneBit bit21(SraOut[21], Shift, DataOperand[21], DataOperand[23]);
    mux2OneBit bit22(SraOut[22], Shift, DataOperand[22], DataOperand[24]);
    mux2OneBit bit23(SraOut[23], Shift, DataOperand[23], DataOperand[25]);
    mux2OneBit bit24(SraOut[24], Shift, DataOperand[24], DataOperand[26]);
    mux2OneBit bit25(SraOut[25], Shift, DataOperand[25], DataOperand[27]);
    mux2OneBit bit26(SraOut[26], Shift, DataOperand[26], DataOperand[28]);
    mux2OneBit bit27(SraOut[27], Shift, DataOperand[27], DataOperand[29]);
    mux2OneBit bit28(SraOut[28], Shift, DataOperand[28], DataOperand[30]);
    mux2OneBit bit29(SraOut[29], Shift, DataOperand[29], DataOperand[31]);
    mux2OneBit bit30(SraOut[30], Shift, DataOperand[30], ones);
    mux2OneBit bit31(SraOut[31], Shift, DataOperand[31], ones);
endmodule

module right_shift_0bit(SraOut, Shift, DataOperand);
    output [31:0] SraOut;
    input Shift;
    input[31:0] DataOperand;
    wire ones;
    assign ones = DataOperand[31];
    mux2OneBit bit0(SraOut[0], Shift, DataOperand[0], DataOperand[1]);
    mux2OneBit bit1(SraOut[1], Shift, DataOperand[1], DataOperand[2]);
    mux2OneBit bit2(SraOut[2], Shift, DataOperand[2], DataOperand[3]);
    mux2OneBit bit3(SraOut[3], Shift, DataOperand[3], DataOperand[4]);
    mux2OneBit bit4(SraOut[4], Shift, DataOperand[4], DataOperand[5]);
    mux2OneBit bit5(SraOut[5], Shift, DataOperand[5], DataOperand[6]);
    mux2OneBit bit6(SraOut[6], Shift, DataOperand[6], DataOperand[7]);
    mux2OneBit bit7(SraOut[7], Shift, DataOperand[7], DataOperand[8]);
    mux2OneBit bit8(SraOut[8], Shift, DataOperand[8], DataOperand[9]);
    mux2OneBit bit9(SraOut[9], Shift, DataOperand[9], DataOperand[10]);
    mux2OneBit bit10(SraOut[10], Shift, DataOperand[10], DataOperand[11]);
    mux2OneBit bit11(SraOut[11], Shift, DataOperand[11], DataOperand[12]);
    mux2OneBit bit12(SraOut[12], Shift, DataOperand[12], DataOperand[13]);
    mux2OneBit bit13(SraOut[13], Shift, DataOperand[13], DataOperand[14]);
    mux2OneBit bit14(SraOut[14], Shift, DataOperand[14], DataOperand[15]);
    mux2OneBit bit15(SraOut[15], Shift, DataOperand[15], DataOperand[16]);
    mux2OneBit bit16(SraOut[16], Shift, DataOperand[16], DataOperand[17]);
    mux2OneBit bit17(SraOut[17], Shift, DataOperand[17], DataOperand[18]);
    mux2OneBit bit18(SraOut[18], Shift, DataOperand[18], DataOperand[19]);
    mux2OneBit bit19(SraOut[19], Shift, DataOperand[19], DataOperand[20]);
    mux2OneBit bit20(SraOut[20], Shift, DataOperand[20], DataOperand[21]);
    mux2OneBit bit21(SraOut[21], Shift, DataOperand[21], DataOperand[22]);
    mux2OneBit bit22(SraOut[22], Shift, DataOperand[22], DataOperand[23]);
    mux2OneBit bit23(SraOut[23], Shift, DataOperand[23], DataOperand[24]);
    mux2OneBit bit24(SraOut[24], Shift, DataOperand[24], DataOperand[25]);
    mux2OneBit bit25(SraOut[25], Shift, DataOperand[25], DataOperand[26]);
    mux2OneBit bit26(SraOut[26], Shift, DataOperand[26], DataOperand[27]);
    mux2OneBit bit27(SraOut[27], Shift, DataOperand[27], DataOperand[28]);
    mux2OneBit bit28(SraOut[28], Shift, DataOperand[28], DataOperand[29]);
    mux2OneBit bit29(SraOut[29], Shift, DataOperand[29], DataOperand[30]);
    mux2OneBit bit30(SraOut[30], Shift, DataOperand[30], DataOperand[31]);
    mux2OneBit bit31(SraOut[31], Shift, DataOperand[31], ones);
endmodule


module right_shifter(SraOut, ShiftAmt, DataOperand);
    input [31:0] DataOperand;
    input[4:0] ShiftAmt;
    output[31:0] SraOut;
    wire [31:0] Bit0Res, Bit1Res, Bit2Res, Bit3Res, Bit4Res;
    right_shift_0bit rightShift0(Bit0Res, ShiftAmt[0], DataOperand);
    right_shift_1bit rightShift1(Bit1Res, ShiftAmt[1], Bit0Res);
    right_shift_2bit rightShift2(Bit2Res, ShiftAmt[2], Bit1Res);
    right_shift_3bit rightShift3(Bit3Res, ShiftAmt[3], Bit2Res);
    right_shift_4bit rightShift4(SraOut, ShiftAmt[4], Bit3Res);
endmodule